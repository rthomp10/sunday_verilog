// **********************************
// Full Adder testbench
// by: Ryan Thompson
// **********************************

module ripple_carry_64bit_tb();
wire signed [63:0] sum;
wire cout;
wire OF;
reg signed [63:0] a;
reg signed [63:0] b;
reg  cin;

ripple_carry_64bit RC0( sum, cout, OF, a, b );

initial begin
    a = 10; b = -20;
#10 a =  5599221927511852972; b =-9073391711843153140;
#10 a =   125843118319673708; b =-7029686126400350234;
#10 a = -6626586882120967886; b = 3892734086233570300;
#10 a = -7567988178298816346; b =-7189453062790077394;
#10 a =   592745535363237000; b =-4295411505309829984;
#10 a =  6778898353225019333; b =-1396929036405534772;
#10 a =   290312938777992501; b =-1693503905809697010;
#10 a =  8575157146419222516; b =-7446083003105828759;
#10 a =  7805619934991066976; b =-2329683517538619121;
#10 a = -8457326708746248500; b = 8933545440415771134;
#10 a = -8384498550222719207; b =-8225720462311965122;
#10 a =  5016413531290329547; b = 1620835055772151393;
#10 a = -2396720075021124139; b = 6565060624351548898;
#10 a =  8756096006914685648; b = 6301982416632616723;
#10 a = -1470614879829494579; b = 7804960753217598729;
#10 a =  8101314306412321434; b = 1696026836459731456;
#10 a =  4547028640344879775; b = 5779657945713253054;
#10 a =   -33533027650960088; b =-8632004510834332950;
#10 a =    23096905326066765; b = 2999616570516881122;
#10 a = -6892050368127303954; b =-7633741690204480755;
#10 a = -6397533401812556077; b =-3133095051764846338;
#10 a =  -983611311585121236; b = 3302033551291320904;
#10 a =  -805828812241324012; b = 4736977790225120819;
#10 a =  1650135588792804994; b =-8419705584332514078;
#10 a = -1904179175795330685; b = 3071518122021549527;
#10 a = -8433565248075562662; b =-4090755593447856424;
#10 a =  -320229163522459137; b = 4466698140372028545;
#10 a = -8365352515154385149; b =-1769744562461170822;
#10 a =  8029209101778457407; b =-1006764421977267873;
#10 a = -7879697700913105533; b = 4349686864040919313;
#10 a = -9178873047882275028; b = 6373368831946348467;
#10 a = -1040351340750794157; b = 6979047705648197226;
#10 a = -7951068199080547545; b =  126450605476960587;
#10 a =   508134022164865434; b =-6778824846222629381;
#10 a =  7445457076962022293; b =  526114371417462296;
#10 a =  7305544011324269284; b = 7582579546691878039;
#10 a =  1541735455966452900; b = 6635438977702751350;
#10 a =  2854214096686148420; b = 8665504473906395854;
#10 a =  -390946583210668124; b =-7330767894173261531;
#10 a = -5952159258982133892; b = 7568652153372798727;
#10 a =  8145744869005091707; b = 4461747306444515747;
#10 a =  5838672863886387925; b =-5767041004222008892;
#10 a =  5960862500006112157; b =-7385299919714859628;
#10 a =  4267292917629836517; b =-6516967423072778865;
#10 a =  4137580239285775024; b =-5149329293057986514;
#10 a =  2643023670507015526; b = 7919885665873411609;
#10 a = -5538938435248079156; b =-3453923133049803546;
#10 a =  8910022516601562726; b = 5594503716843436989;
#10 a =  6909142613382597738; b =-1218515048110619699;
#10 a = -2386127518659592150; b =-6846767655301744517;
#10 a = -6815849060657679249; b =-1228202050904613620;
#10 a =  5714779459212850260; b = 7190423059372391560;
#10 a = -7255729558549911617; b = 7987520561947225693;
#10 a =   948429068982750254; b = 4005140714472405259;
#10 a =  7796570658536682580; b = 6990487115605157645;
#10 a =  -637888390100998310; b =-3077813523392619824;
#10 a =  4238264959324070591; b =  -37965819277855933;
#10 a =  6269537513499946930; b = 4134729987642894407;
#10 a =  8834074481322271560; b =-3518289805054397606;
#10 a = -6310058247795273022; b = 3512022914817055364;
#10 a =  7289839610128698002; b = 4762495609653693642;
#10 a = -5766864379392692915; b = 5553070326130275748;
#10 a =  8338095794085366770; b =-5954190803751878943;
#10 a = -6687412454855600462; b =-8619334172319419082;
#10 a =  3893242104366499047; b =-9165869667202848176;
#10 a =  8719075204911463153; b =-8507833250647803401;
#10 a = -7926563180461026709; b =-1317678225756220373;
#10 a =  8530703474273415522; b = 8886787539172512471;
#10 a =  -707292090388796837; b = -597562586826919610;
#10 a = -5568953431868867803; b =-4278512197784715079;
#10 a =  7162696349164539316; b =-8616280970915535594;
#10 a =  2262954627082897455; b = -952108641040262449;
#10 a =  9163926912051408919; b =-5587910976516935099;
#10 a = -1039504208308413341; b =-3484959141908494153;
#10 a = -1291381655351215929; b =-7010161366924896408;
#10 a = -7904793985155824385; b =-5050153574774556194;
#10 a =  4006160316257963978; b =-8222299613140769351;
#10 a = -7446065508060833246; b =-6309413587358137169;
#10 a =  1262419794867128548; b =-4276614964675721420;
#10 a =  1751456881694440961; b =-7274339214520866937;
#10 a = -4085388555879664056; b = 8450845718521114532;
#10 a =  4216248319607783962; b =-7590471841133101065;
#10 a =  8533299366624320697; b = 8027181867091708274;
#10 a =  6576697536743217414; b = 6545933559562767488;
#10 a =  6781426785887839639; b =  238407136350082993;
#10 a = -2693901759088158434; b =-6577229211369974689;
#10 a =  -211816726161178383; b =-4416046730106523072;
#10 a =   744057974788159557; b = 3220675450320581175;
#10 a =  9015983165379053728; b = 2112882073917560644;
#10 a = -8158065906043417836; b =-1789069408030687465;
#10 a =   383055310195961177; b = -495070620188503203;
#10 a =  7687556311610769876; b =  -77202853514632489;
#10 a =  -112403483484376159; b =-6426219444353793776;
#10 a = -2726192894151558144; b = 3633604397126517419;
#10 a =  2432248309655379617; b = 1462387551669124485;
#10 a =  8117086711331535833; b =-7220054846226708130;
#10 a = -2315347405599032881; b =-5867863910359211558;
#10 a =  2825914046407054633; b = 1851752032326851072;
#10 a = -6237299360291849304; b = 3905821927579375032;
#10 a =  2333485990445799260; b =-9044627570319684964;
#10 a =  1799919859778032655; b =-8891923922670447178;
#10 a = -2457246499902826170; b = 3985259948272440346;
#10 a =   818893172777320831; b = 2423818169767853827;
#10 a =   864337286297994358; b =-8091068663498576611;
#10 a =  8531051160075798563; b =-6385772176720385167;
#10 a = -1409713208221841321; b = 7617093056574369491;
#10 a = -4017138349483852795; b =-8939599338766473322;
#10 a = -8853505449226503787; b = 2206515053695753064;
#10 a =  4314494103137216457; b = -725645920376201718;
#10 a =  5540353769901191608; b = 6358677148316200253;
#10 a = -5016909398242867218; b =-5009839040939351244;
#10 a =  8345881517115067506; b =  382607450714723168;
#10 a =  -574995337915262947; b =-3842926097570983191;
#10 a = -3489893239915534920; b = 8648681654181034987;
#10 a =  6471176958025481306; b = 6084824854556974980;
#10 a =  -425887340308326840; b = 6942707179982807808;
#10 a = -8662111769287919167; b =-8749096620928333422;
#10 a = -6988264116314976835; b =-1985958544537700829;
#10 a =  6129909720897268353; b = 6633833414352924018;
#10 a =  6723550814019034978; b = 2950654430716185580;
#10 a =  6647510423368806373; b = 5704442870987262752;
#10 a =   282544591555605642; b =-8304547994470863468;
#10 a =  7528067868072734529; b = 4395966877659760915;
#10 a =  5351247057272803721; b = -219499273512881426;
#10 a = -6919532060470875258; b = 6508602873738272140;
#10 a =  2917149809422391764; b = 9204470314989965397;
#10 a = -3137091962089575286; b = 6855016823129791554;
#10 a =  -246851826206799052; b = 7406543434817331687;
#10 a = -2621267972981203723; b = 4951573665182363644;
#10 a = -6067115272846651878; b = 6982102946174737878;
#10 a = -8060366874062312540; b = -688729053275174085;
#10 a = -5628079961872236166; b = 8825923690017524054;
#10 a =  1599943223397786290; b =-7889044043089268377;
#10 a = -5636400626460622924; b = 1943243305826297075;
#10 a = -3371569370708916184; b = 1179285147392821846;
#10 a = -4363746415012493924; b =-2029622618012604500;
#10 a =  1788383771996546784; b = 6675982753196639811;
#10 a = -1982591943019212063; b =-8787550022613560008;
#10 a =  -890218766641702809; b = 5257832702547293605;
#10 a =  5785181496982417827; b = 6040815099718229315;
#10 a =  4781888999353752466; b = 6274118193166079596;
#10 a =  7673540953670151460; b =  163143140257471818;
#10 a =  3094555051400740999; b = 1637477871578921269;
#10 a = -5048695002948525464; b =-4281969165932202460;
#10 a =  5237619560122580601; b =-4098410925661316177;
#10 a =   182508943049381754; b = 4203008557973051743;
#10 a = -2710605822329480426; b =-5978608711670002161;
#10 a = -2296680730491138245; b = -758564511049818350;
#10 a = -8816771296227887846; b = 3476698358387008402;
#10 a = -7967804632574327792; b = 4086576009279640399;
#10 a = -1923555456168791393; b = 8846689731725571393;
#10 a =  -509491550915713990; b = 8544246629349879867;
#10 a =  4194115558563370138; b =-6742202317196833755;
#10 a =  1455044463595001978; b =-1495184219704327859;
#10 a = -7138637764571973903; b = 2141129573436380672;
#10 a =  4735427883456944171; b = 6807492117484349989;
#10 a = -8297276190861705157; b = 4076463507034792240;
#10 a = -2037385669166870472; b = 3351109022536281670;
#10 a =  2790132534028478860; b =-1702349955069379335;
#10 a = -5948594702426347711; b = -260832556842157694;
#10 a =  3341695706333251304; b =-9216927306675395285;
#10 a =  4728183419013217065; b = 6731341437260808712;
#10 a =  1596887168224310089; b =  417689964541207257;
#10 a =  1413762954249691536; b =-1296312289413111576;
#10 a =  7211944393904702811; b =-7313590257225140129;
#10 a = -5921268540210684752; b =-7988678388620043920;
#10 a = -7495773448130646194; b = 5070773443877614773;
#10 a =  8414732564759594875; b = 6589498388047073932;
#10 a =  7394967475613721218; b = 1068444613920370015;
#10 a =  2408473284348918729; b =-4518654658461767742;
#10 a =  1648559816137469443; b = 7016057952031012781;
#10 a = -6199949358767468112; b =-4924405635496226076;
#10 a =  3502469614332576126; b =-7150913321770824925;
#10 a = -5562961411668983946; b =-8171161551368829980;
#10 a = -2208921609778702394; b = 1595006087527818717;
#10 a =  4070671681169862944; b = 6416702717914218342;
#10 a = -6890838674334252191; b =-1155434380248455822;
#10 a = -6504487425048985538; b = -644014037852099286;
#10 a =  4431665120158562905; b = 8538197010630021276;
#10 a =  6006623468393946058; b =-2718769740776834386;
#10 a =  4765885012792048290; b = 4586421410478029658;
#10 a = -7829917923791059488; b =-7107771688129375490;
#10 a = -5595186958130495050; b = 1113280797883520053;
#10 a = -2175590252804086415; b = -240259237043473239;
#10 a = -2412541986440881078; b = 7698595875410516944;
#10 a =  -741035488564604095; b = 4518299650332825769;
#10 a = -7793450099634144433; b =-4042945654761763063;
#10 a =  4865609926133095086; b = 2873208530239942819;
#10 a = -3145954933537851437; b =-5615829776132582096;
#10 a =   -63566772783624883; b = 7109568255813754581;
#10 a =  -178261978143301967; b = 2566759521676904779;
#10 a = -5354933876210937023; b = -714590249916822915;
#10 a =  2583868074628639716; b =-3240866649601670320;
#10 a =  7701850048359035232; b = 3670708648649768222;
#10 a =  1909412735828891252; b =-8958816258008897136;
#10 a =  2015669775480937234; b =-4230617939863287182;
#10 a = -4254275357477779809; b =-9093672534700133031;
#10 a = -3126725999879102504; b = 6077252973351313399;
#10 a = -1895382705383207879; b =  569707070885383544;
#10 a =  1901384613167011887; b = 8273248178331175696;
#10 a =  2078948419885665532; b = 5502859595967247290;
#10 a =  1097965373362184150; b =-2304855382315205505;
#10 a =  -998525441645594862; b =-8509328755271450056;
#10 a =  6695841463746080255; b = 3538674199257254711;
#10 a = -5159076378039626734; b = -272284914038094262;
#10 a =   290394676418383645; b =-4683550479335858849;
#10 a =  6706719726660604199; b = 3961439101092508553;
#10 a =  5875027599019537277; b =-7548860498939323475;
#10 a = -7953007242656803656; b = 5199103333983582175;
#10 a =  3598286275300261956; b = 3294845053905274865;
#10 a =  6451676350548604088; b =-9146635523445992318;
#10 a =  -880702070047010949; b =-7442968733763892365;
#10 a =  4431787183339578448; b =-1646665860596597973;
#10 a = -3266714066946699053; b = 4882901422412927603;
#10 a = -5441517265935394240; b =-7872867665755229334;
#10 a =  7211392450993342519; b =-5913598157519829054;
#10 a =  4138981247468602798; b =-4732104960610158098;
#10 a =  4049315762301466853; b =-8161200399650065646;
#10 a = -6965468699193858847; b = 6717711416395867084;
#10 a =  7940030719377733418; b =-3546931943693176003;
#10 a =  4337445661893136742; b =-2451511040730532571;
#10 a = -6523011041163790357; b = 7761249482825822941;
#10 a =  1165964451569980013; b = 5857305876658829383;
#10 a = -2843511997966350343; b =-4564865506242560492;
#10 a =  8656410509924073908; b = 4402593517146070357;
#10 a =  2530206813867962791; b =-4146237617254441870;
#10 a = -1117101610790619958; b =  341900831991869079;
#10 a =  4626561213614103103; b = 1242976384763903396;
#10 a =  2974683091453563480; b =-8116124587107899124;
#10 a =  4947001522910468656; b = 5602408392374931448;
#10 a = -7909690184094452107; b =-6753292157131616878;
#10 a = -6264886440499460914; b = -739258824522604249;
#10 a = -6825475857035840592; b = 3378416711909031699;
#10 a = -3510263970520730670; b =-3083008843629961452;
#10 a =  4897616711797245664; b = 1412923286305860952;
#10 a =  7047202071394582657; b =-5100328138027348799;
#10 a = -4258543309232370315; b =-9128916352179013458;
#10 a = -2765367946413424638; b = 8880253541292040179;
#10 a =  3108506991900733480; b =-7689159359259788749;
#10 a =  8625647422428801919; b =-3051780755122893799;
#10 a = -6649432747536646420; b = 6869005756576849628;
#10 a =   224959883787664456; b = 6467879041020026539;
#10 a =  3696485514032648573; b = 3276564577355576537;
#10 a = -6518000392526563322; b =-7266795968470231618;
#10 a =  6998930740635559494; b = -803823134850649054;
#10 a = -4169740089997849140; b = 8798068332628252986;
#10 a =  7517504532195213650; b =-7660985760923005344;
#10 a = -8431716696716516752; b = 6149518764919839651;
#10 a =  1473498067362439700; b = -641644037964145122;
#10 a = -2468259106858029046; b =-7270012361669310844;
#10 a =  6689940896216870353; b =   57522910861383843;
#10 a = -5086654316291101284; b = 7397188741628329166;
#10 a = -5162115080518915325; b =-6739004664949510863;
#10 a =  6515908336312600121; b =-7422902436291887715;
#10 a =  1823197532519013516; b =-2756917895112997917;
#10 a =  6483782794833817541; b = 8066978003439092934;
#10 a = -3388098624345258763; b =-3476071623891561054;
#10 a = -3399639883882977487; b =-7241044537356437674;
#10 a = -4632413741034752774; b =-5380476081503390335;
#10 a =  5101125258080915380; b = 7024717838588121557;
#10 a =  7011918523199095484; b = 7674499487637461731;
#10 a =  2587968398052847487; b =-3518478093577667209;
#10 a =  5202751479003169140; b = 4482725693650481394;
#10 a =  -555876413379425090; b =-6404665476963851884;
#10 a =  4264417508385920525; b = 6565129862207554876;
#10 a =  7639731349228030042; b = 3088067349986100518;
#10 a = -2554534591973320728; b =-7512126165663220999;
#10 a = -4960945430234056348; b =-7461789457350517220;
#10 a = -4301535952856451070; b =-8746250600816671283;
#10 a =  8276778903586540135; b = -469669146872767858;
#10 a =   979494924224180082; b =-8762124820975865097;
#10 a = -3363969026379459270; b = 9170571801518263899;
#10 a = -5710554188179142668; b =-4694447095105650722;
#10 a =  2500815882078454725; b = 3508107426242290112;
#10 a = -1693021614498396234; b = 4127947155606249567;
#10 a =   284722250467243531; b =-1187724609641278347;
#10 a = -5737963953210277314; b = 4404677667367190707;
#10 a = -8495260404578939880; b = -611984082207096242;
#10 a =  4163737213853092044; b =-7738581286562995096;
#10 a = -8463977919119608565; b =  216796824212704180;
#10 a =  4420359639715072678; b =-5874662724873159487;
#10 a = -4598191881274330212; b =  485587508377657779;
#10 a =  5870042728044797946; b = -597870544276487523;
#10 a =  5299670305864028521; b =  376696898269440519;
#10 a = -8405968114169695962; b = -404918199411203581;
#10 a =  4213102989492704099; b =-7354248716658342552;
#10 a = -6614763913445302523; b =-6958727530642085071;
#10 a =  3632295591674555849; b = 1012094061912485933;
#10 a = -3646967100891944736; b = 3610202679540587350;
#10 a =   295722438467388314; b =-7511846009542652541;
#10 a =  4111254361244212126; b = -942367885739980224;
#10 a =  6982994341542183893; b =-1617015717841755361;
#10 a = -5363995474213189266; b = 2496542212558817797;
#10 a = -9112200299893404016; b = 3715214068057247268;
#10 a = -4484487234594872969; b =-8554788624537489607;
#10 a =  5392485228544547718; b = 6552883489187762061;
#10 a =  8099857894663327332; b =-5196863392934474715;
#10 a =  9117268882788977419; b = 7899795439629296349;
#10 a =  -541886820470639245; b =-4763796954911646716;
#10 a = -4627982329972192767; b = 7596786472334334172;
#10 a =  1898346180168102682; b =-7041550908479863884;
#10 a =  5561482709590100662; b = -620644778872560535;
#10 a =  -215746691760331595; b =-6451946800005979003;
#10 a = -6135972907417130732; b =-1418831750100288792;
#10 a =  2379806969749322970; b = 5764712034986529812;
#10 a = -3498751230870494020; b =-6939607465901944448;
#10 a = -1487455866814883264; b =-8804575747845586754;
#10 a =  8617176780018446178; b =-7458869898515218377;
#10 a = -2350018545849529271; b =-6452464650274626618;
#10 a =  4706359959592454572; b = -777199251347083795;
#10 a = -3071436730142217488; b =-5607587302102483415;
#10 a =  6367682836845236258; b =-8591848888615321236;
#10 a =  8555635846237030596; b =  -62497717879514791;
#10 a =   141732845137224200; b = 2634853653436192683;
#10 a =  7355656986968375131; b =-4093378952795192961;
#10 a = -2206841416270030300; b =-4279929385962734864;
#10 a =  1596039600969390471; b =-4230865085780046340;
#10 a = -6260444103224374637; b = -697283190479987600;
#10 a = -4138012997039283930; b =-3144648556565398668;
#10 a =  8735055330761243594; b = -885933351550445909;
#10 a = -7858848940922788358; b = 7920588674543631875;
#10 a =  -825042847919412677; b = 8424080224136447125;
#10 a =  4036894687723632795; b = 7528664361327287530;
#10 a = -7958084347552686295; b = 9221443684601711717;
#10 a =  3235606384811158131; b =-2193150426281934286;
#10 a = -7021703128777896832; b =-2641747589790126505;
#10 a =  4660113176761783672; b = 5401317844103077650;
#10 a =  7163808051786654507; b = 4374339502590793909;
#10 a = -1792655772650128963; b =  298566485876682853;
#10 a =  7376244146389157350; b =-2237678228809674469;
#10 a = -5733446417664310283; b =-4867676910915670274;
#10 a =    -3220151069313831; b =-1242344540040682379;
#10 a = -6829958027245605925; b =-1461866193287798246;
#10 a =  1717466935558921910; b = 3570108677077047780;
#10 a = -3999334021550608789; b =  719443786059269025;
#10 a =   818423751062414101; b =-5438387959171568895;
#10 a = -6689991455350785774; b =-3115311363921168323;
#10 a = -2981042845393057916; b = 2916507841259570291;
#10 a = -7720513342334978748; b =-8581753677496976320;
#10 a = -2230505630210113588; b =-5002545803414941972;
#10 a = -3991230454239236425; b = 3753910579860683844;
#10 a =  -576339937844889249; b = 1047731815806606920;
#10 a = -8195703849722245666; b = 5890707721768228764;
#10 a =  -982049056853925308; b =  907610892740145962;
#10 a =  7722878645745107645; b =-5670761424140884162;
#10 a = -6999394452190968804; b = 9017276320639811633;
#10 a = -8129507479482311003; b =-3605096774474202045;
#10 a =  5919821213505832710; b =-6143471463296422585;
#10 a = -3829826906296816371; b = 4727920265476985621;
#10 a = -3386652710402951212; b = 6692990013381983681;
#10 a =  7514981863214040793; b = 5279406596077159285;
#10 a = -3580964522476445932; b = 4485447781733713522;
#10 a =  7558550074027701365; b =-3945158878798175412;
#10 a =  3022896743049559707; b =-1737196216955589090;
#10 a = -8056698518455676448; b =-1813840610518877195;
#10 a = -1548040941394349467; b = 6190053941970433855;
#10 a =  8645689108882077238; b =-2801330880423410441;
#10 a = -4826489842529374112; b =  894776075583214047;
#10 a = -7880395837333524092; b = 2482851747316267168;
#10 a =  5960133500518213229; b = 5626755216979156886;
#10 a = -3484464729632447872; b = 3372575080638040673;
#10 a = -3022123879835407776; b =-2396091772178868706;
#10 a =  1969142091711213484; b =-3599182826107316875;
#10 a = -8745470179216043008; b = 4249530689550941892;
#10 a = -1976784043695059721; b =-5637280014353627062;
#10 a =   889113550945730012; b = 2817385673582448694;
#10 a =   412287001603402695; b = 5938896371340281283;
#10 a =  8901407120933776971; b = 7992513418240635414;
#10 a =  4712811152317364063; b =-3555626937785447084;
#10 a =   954974931834428099; b = 5859459762679823680;
#10 a = -6173254902049145975; b =-7501241334519795014;
#10 a =   563066685582752495; b =-7506406955054502553;
#10 a = -8340630454775687239; b = 5727220616620431154;
#10 a =  6860732178871975555; b =-5740363575988539443;
#10 a =  -610899172384038191; b =-8690641286213023900;
#10 a = -1701853478155814260; b = 3068628693436731632;
#10 a =   -84894192107665077; b = -179287416467468002;
#10 a = -1695865776263885239; b = 6832675962310918536;
#10 a =    91481830147367287; b = 5036664163826101661;
#10 a = -6745787169388071482; b = 2356566511331855716;
#10 a =  5416155468854556487; b = 8063041005143554663;
#10 a =  6313246495093008573; b = 3460209990654375833;
#10 a = -7606542739318825753; b = 5437546286373431722;
#10 a =  5284554888064558975; b =-6069711902037440515;
#10 a =  -798659265678465474; b = 8040455165469802533;
#10 a = -5360462105843226919; b =-6928449929309673277;
#10 a = -1543758523880702319; b = 7358751126517832168;
#10 a =  1277060530670171332; b =-3518961839302465863;
#10 a =  8184364170550415897; b = 1949498605757725807;
#10 a =  1904813634680841672; b = 7334452814980077996;
#10 a =  5166065496237290772; b =-5584167211071591744;
#10 a =  4359478271445217674; b = 5575921050192964241;
#10 a =  -124659716738108069; b = 8714282176631777025;
#10 a = -8185384531911144583; b =-6644401005421874629;
#10 a =  7433751246498984379; b = 6628025103305420360;
#10 a =  8882217496154189536; b = 5781499921168007250;
#10 a =  6123264568455102147; b =-2936238653158603251;
#10 a = -1133211782803976416; b = 2469261358762748507;
#10 a = -3639320281453875406; b = 2678034872002694318;
#10 a =   592776260151197411; b = -880725918650895356;
#10 a =  3988347153438340227; b = 7669412702740987786;
#10 a = -3161354467980521751; b = -176358541252829381;
#10 a =  5385322412066173554; b = 5952322865178819648;
#10 a =  3886077837972469192; b =-4049017109616524896;
#10 a =  5991532003682335914; b = 2280380539206700158;
#10 a = -3846158735321673061; b =-6084492576291316218;
#10 a = -3868555578708114558; b =-7119506608604134837;
#10 a =  1683666999029314666; b =-4646814812368182640;
#10 a =  8376415113683347187; b =  410662861018152338;
#10 a =  4527538211488810872; b = 4867818914292215315;
#10 a = -4895929609266201490; b =-2415431481454357026;
#10 a =     1693699535246450; b = 2592068319346176028;
#10 a = -1229274940893594235; b =-1662094639115539936;
#10 a = -6728731084523562236; b = 9166889820989869896;
#10 a = -3889487079876498519; b =-5770518389216234904;
#10 a = -1514731060224110352; b = 7845398570224913798;
#10 a = -5209981776514334032; b =  289544814333286365;
#10 a =  2493767907273644575; b = 1474201881231939762;
#10 a = -8942099268628464378; b = 2779023112249001473;
#10 a = -5345934932825767167; b = 5530371213844265539;
#10 a = -2339233383827529246; b = 6794293985413881622;
#10 a =  4603587033248998890; b = 5814159878525816488;
#10 a =  7257504124655091032; b =-1750423620919040499;
#10 a =  1570161686032190129; b = 8621790199592082648;
#10 a = -4808573067386457285; b =-6863299988282644593;
#10 a = -7688553525641375281; b =-3343170553859491866;
#10 a =   189872427595545610; b =-6680060936016598203;
#10 a =  -995808632283933115; b =-8425952962648491201;
#10 a =  4480954528899013829; b =-2263560820744265371;
#10 a = -7014243668706503121; b =-7464947393735822558;
#10 a = -3979441021631235843; b =-4753639408897939141;
#10 a =  1358066160571106074; b = 7080719011134467365;
#10 a = -2203154204253109537; b =-3712245809697508127;
#10 a =  8947691589359780842; b =-5824998587880568917;
#10 a =  4391874205305910395; b =-1615433545411631410;
#10 a = -1138266230072755834; b = 2825231209549028012;
#10 a =   661955298355112168; b =-4830615096760899213;
#10 a = -7288236513438889108; b =  737363299159159152;
#10 a = -4512903439851010055; b = 6746979396664203120;
#10 a =  -692808210133112751; b =-5648238319529619026;
#10 a = -1564226404175500759; b =-2137933877817360124;
#10 a = -3488769138840075815; b = 6461497195369022190;
#10 a = -6151102471751249212; b = 8249400811125843863;
#10 a = -3524282682236397895; b =-8386208015766122668;
#10 a =  6563810136954956811; b = 7371346632354525125;
#10 a =  5524968048874725502; b =-6138917491405110754;
#10 a =  3975856565559273950; b =-5992058124406342804;
#10 a =  8214825206680363582; b =-4888937578628604130;
#10 a =  1878251557392532820; b =-4612172507655481528;
#10 a = -7201737568098153472; b = 7111665018708611334;
#10 a = -3223121534626487861; b =-1524249642225466243;
#10 a = -5415759519763764191; b = 3095071087365788415;
#10 a = -4265988069140113008; b =-3345065206133952989;
#10 a =  8276108618132405614; b =-6343653278027117901;
#10 a = -5641027037525385471; b = 1822952017121547915;
#10 a =  8092365071540245480; b =  772033328963151598;
#10 a =  8581654588294005670; b =-3098649179751373870;
#10 a =  -865434773076714488; b = 5887888527934573241;
#10 a =  5592724197477283979; b =-4705418737982665848;
#10 a =  6748624485613505136; b =-3474146700488883248;
#10 a = -4531019998303493037; b =-4711822263274979168;
#10 a = -8534554223159583368; b =-4078449822150738570;
#10 a = -1957444654085462646; b = 6567761361755393525;
#10 a =  7067137442952525069; b = -424369441213167372;
#10 a =  5944546398103501670; b = 7491332230169835883;
#10 a =  6499302309653577795; b =-5044107452804654176;
#10 a =  7495952821728919633; b =-6080832874929208233;
#10 a = -6411571323225330956; b =-8246392628291634494;
#10 a = -4698854580796199338; b =-4270072492385980289;
#10 a = -9095346695035368823; b = 8870740054590063519;
#10 a = -4531425993504545890; b =  240904992087171914;
#10 a =  7072127362119517810; b =-8332736686755500322;
#10 a =  5811925829962314792; b =-1239827082118983401;
#10 a =  5919427321198869569; b =  419169273917803596;
#10 a =   348547945368087676; b = 1888001166017155668;
#10 a = -1757648815611350654; b = 2125031615349850681;
#10 a = -5918002076084756933; b =-8635252003092349122;
#10 a = -4160980775321712625; b = 6325367039931931928;
#10 a = -1828193085527935540; b = 4516257473545318289;
#10 a = -4681181869032284890; b =-2636554913197238456;
#10 a = -5083121754590127405; b = 2627019985135217774;
#10 a = -4831655628877321065; b = 2313401121370814482;
#10 a =  6868534480839981100; b =-1261346118734783115;
#10 a =  1042077087850022967; b =-5036204683284610732;
#10 a =  4783043681111874020; b = 5506280524662143039;
#10 a =  4139072039477881929; b = 1436497608527055564;
#10 a = -8976001629291010126; b = 4567411590596689105;
#10 a = -5163059892323358772; b = 1901579768826282663;
#10 a =  3883249843134684954; b =-2986197199569489110;
#10 a = -8935550112378791685; b = 1743584409442195831;
#10 a =  -344412357021841709; b =-7047718004204535997;
#10 a =   909852276851739079; b =-2906829423892651127;
#10 a = -8170865470582247684; b = 9198140724155674064;
#10 a = -6340391807891757618; b =-2286053149935796329;
#10 a = -5412716942372318160; b =-8608975328090578135;
#10 a =  6564109048861754582; b =-9030939783989545603;
#10 a =  6153163862389609426; b = 7247344062853081366;
#10 a =  3303398178079105145; b =-5501846869422165485;
#10 a = -2499939993452686332; b = -961590516125075805;
#10 a =  -328934335107614854; b =-4160267154943738819;
#10 a = -2578813702118459377; b = 2791308242917927957;
#10 a = -8848694990896560352; b = 1768797097015433691;
#10 a = -3183222641446598564; b = 1499372749352757073;
#10 a = -2822479541875211651; b =-5650292216747161761;
#10 a =  6830903736211777776; b = 5985060924929808137;
#10 a = -6090075290508076478; b =-2083848231505012583;
#10 a =  -331471758952360634; b =-8110268276411372846;
#10 a =  8953293621394402407; b =-5834578442990062287;
#10 a = -1863756299374050949; b = 7821426229610478699;
#10 a = -2363546669590459336; b = 7098498696608486761;
#10 a =   669995587174379069; b =-2195717928453241958;
#10 a =  9113457830955203377; b =-2446967230008331694;
#10 a = -6929964557134983413; b =-4208682711966007422;
#10 a = -3120656792135646239; b =-2181899788214118383;
#10 a =  4641218644065326076; b = 3126171402917798206;
#10 a = -1194120614558441217; b = 3856218335190828472;
#10 a = -8911677222412596900; b =-8684357737432157130;
#10 a =  6669970890662570793; b = 7999120278838197656;
#10 a = -4123243103361631154; b =-2172655084164405615;
#10 a =  6809734625022900656; b = 5686559603597943888;
#10 a =  8646249654095314554; b =-1753174893759818064;
#10 a = -2620829779312040505; b = 1219755350032322263;
#10 a =  5549031456025379457; b = 5637382020653599906;
#10 a = -7307953418617462931; b = 6191851304259271954;
#10 a =  -158942599283220664; b =-5782884182214910145;
#10 a =  8674634017346028750; b = 8938362499436055433;
#10 a =  3593996915835667055; b = 3416091258824166732;
#10 a =   327513992924917154; b = 7178639057409954555;
#10 a =  -723974637181568477; b =-5491760098277317301;
#10 a =  6292583692144083408; b = 2942615312400527717;
#10 a =  4807917365437665061; b = 2594950730328247234;
#10 a =  4096754844317924001; b =-5833697724306841793;
#10 a =  -839288586196831545; b = 3231085994501720683;
#10 a = -8240296480935904563; b = -115291235171280507;
#10 a =  -650347853225236378; b =-1251727866817085058;
#10 a =  8091285149239068006; b = 2489791947318280742;
#10 a =  8413568011923058603; b =-2504741617389496377;
#10 a = -3356525558748144082; b = 3488294172973297647;
#10 a =  4331216103208915539; b =-4777297480217461793;
#10 a = -9178579073164851712; b = 5589711748847307847;
#10 a = -7035734307538135191; b = 1604158165949599997;
#10 a =  6459929100038585682; b =-7343039097780215511;
#10 a =  4304498933459073413; b =    6997806394006572;
#10 a =  8011060326434184096; b =-7007373322657596118;
#10 a =  -149968111974628319; b = 5656660961784272588;
#10 a =  4034162666294108634; b = -588159868884999281;
#10 a = -6340906917976228487; b =-6074242099699495548;
#10 a = -5656165569999374638; b = 8254635549959090921;
#10 a = -7026576379918423015; b = 8993436803488274546;
#10 a =  8493886159588140836; b = 8753089368433458563;
#10 a =  6555949487326478520; b =  593078217709202067;
#10 a =  1801970937331642652; b = 3897563671539843950;
#10 a =   857065949864415653; b =-3740051360959467540;
#10 a =  8040523269034624782; b = 1216996793789582852;
#10 a = -2110820555563298408; b = 3134389354908589215;
#10 a = -6780316773731684271; b = 1854186173347324448;
#10 a = -5321622550743063567; b = -900652589373201000;
#10 a =  8317478680549628802; b =-4869682116258030005;
#10 a =  4585056589967931512; b =-1698127403801271028;
#10 a = -4776230033175477615; b = 5095964021964683241;
#10 a = -8469913670993418689; b =-3347902451371233885;
#10 a =  5350407008264303272; b =-2471683660182143677;
#10 a = -6765112617475304941; b = 5062088773604603011;
#10 a = -6034977774239197206; b =   -2639112711632208;
#10 a = -3712169382773618294; b = 1702473287114919553;
#10 a = -8705043045874496624; b = 6249105084425509726;
#10 a =  5029553776964783071; b =-8205637755288531206;
#10 a =  2293458359368605186; b =-6664193977457024723;
#10 a = -6513687724396847034; b = -362915899597588943;
#10 a = -2301773253335438673; b = 8765362993559799161;
#10 a =   135947485410855383; b = 1275296518166572638;
#10 a =  3917825424262420502; b = -729205852476211496;
#10 a = -3385661109695336833; b = 6666156466775539635;
#10 a = -6340820627065720910; b =-4284361819171812308;
#10 a =  6654634507970439917; b = 8631652466949945940;
#10 a =   -86351464684370003; b = 7861354887795000990;
#10 a = -8284282770155792821; b =-1340762047962426534;
#10 a =  5943888392098911928; b = 1740236369849302932;
#10 a =  6933423141572184943; b =  184254854261519596;
#10 a =  2333977918171061849; b =-8747985733692284132;
#10 a =  8305828801596010199; b = 8096061443495553436;
#10 a =  9042245854639754478; b =-3274263351986865990;
#10 a = -4715421500133149446; b = 8512483160977618295;
#10 a = -6457176759075702768; b = 6596369584065467273;
#10 a =  8343803439961333529; b =-5975384429774817412;
#10 a =  5534355883401750448; b =-4860596902790086424;
#10 a =  3258454872337022366; b =-5757232476640913770;
#10 a = -6922040805390544352; b = 5713574058932965123;
#10 a = -6315091746620141553; b = 2499321051830178810;
#10 a =  2146763252199275954; b = 3871655627417008328;
#10 a = -4061734593845697619; b =-7838753381608649011;
#10 a =  3852314424523806204; b =-1893392696541270642;
#10 a = -3902751588670726226; b =-6062978886660471067;
#10 a = -8817654179804298061; b = -972126085265179216;
#10 a =  2000299678933242651; b =-6687018654465702244;
#10 a = -3798880384891508555; b =-5532160491044192912;
#10 a =  3191574271727039250; b =  864100556004810739;
#10 a = -2542476092908840955; b = 4926483438617010151;
#10 a = -8871567547332352816; b = 7010047985412161805;
#10 a =  8845444003561321934; b =-6461968513746270283;
#10 a =  8681010436700977392; b =-3933114469920703293;
#10 a =  3818010063915537639; b = 2059071460825229897;
#10 a = -1806269656066725163; b =-8234226342242216102;
#10 a =  6445283910246707729; b =-3138930546637042650;
#10 a =  9009238830759681473; b =-4807021844631389605;
#10 a = -1772720584286786964; b = 3355628044428102056;
#10 a =  8693563406365109188; b = 4149663763804149398;
#10 a =  6250472244265097267; b = 1194649068495695476;
#10 a = -5582791041528451758; b =-2635613830828753856;
#10 a =  1286478731646223615; b = 8920318044565443645;
#10 a = -2335898648626891640; b =-7826363312097294697;
#10 a = -4703699012331208901; b = 1022634130463850067;
#10 a =   221526320613347490; b =-9068627997701073716;
#10 a =  2603527876463420386; b = 8109938576013563985;
#10 a =  8225300361993749201; b =  405514086961075691;
#10 a =  5407412202484855434; b = 1933164654681877958;
#10 a =  7427684284140729446; b =-4300087896137491300;
#10 a =  7617085063097743606; b =  871534725409330443;
#10 a = -7478447821666815238; b =-7826313382928752706;
#10 a =  5648435409514275112; b =-1920205535735052103;
#10 a =  5269135444342655978; b = 7744325911378861079;
#10 a =  3665308967997541376; b =-3578590856070603147;
#10 a = -6479876818575529269; b =-5571630390481619666;
#10 a =  8913639656173103861; b = 2244272928880637597;
#10 a = -2914981038679492868; b =-5564586901792628320;
#10 a =  2824836913380102004; b =-8766103540212792541;
#10 a =  5846533573578583676; b = 7116286164904294061;
#10 a = -3774459894354766662; b =  264417132352853433;
#10 a =  8085127689142036541; b =-4783469383099744581;
#10 a =  3225388113534785790; b =-8010403725877540074;
#10 a = -5645126874504086412; b = 3213624543324013716;
#10 a =  4394434453492035424; b = 4596548051728315586;
#10 a = -8442395293608344882; b =-3142495062333665225;
#10 a =  2040424608467966505; b =-3745754111944943798;
#10 a =  2403629153284792244; b = 6600871991585721262;
#10 a =  5620813261852069259; b =-8303484699326957042;
#10 a = -8184203259125156293; b =-2399741994988206622;
#10 a =   476775499910913108; b =-4846641676243033159;
#10 a =  3911866649975020205; b =-4328617366739886365;
#10 a = -7543430739877304140; b =-8110289564049020836;
#10 a =  7280298915361220247; b =-6310932202178438549;
#10 a = -4859863070465728110; b =-1384607991727521113;
#10 a = -1264075689235889881; b = 6171494587219062478;
#10 a = -3276752213009503362; b =-8702692812734026549;
#10 a = -3865835064182025911; b = 8924031334902435178;
#10 a = -7947014772879094944; b =-2083260657773301920;
#10 a = -2530726748016649626; b =-3344913852617892116;
#10 a = -6072325146991891271; b = 7344062752447046999;
#10 a = -1881828615779527153; b =-2698362937042404585;
#10 a =  -818569030924571564; b =  664090329916573620;
#10 a =  3546696543644757031; b = 1004762216856333793;
#10 a =  -955806320459699922; b = 2998773216155370727;
#10 a =  8667870030772866796; b =-6176622140420521889;
#10 a = -3002596817949790218; b =-6512074220689322678;
#10 a =  4673445873018820137; b =-3563246541747050128;
#10 a = -4256276977054378131; b =-2683592657606895160;
#10 a = -2627796886901723676; b =-3931799913425672386;
#10 a = -8883301795551580386; b = -892094303574161406;
#10 a =   671193082135255278; b =-1831724870521664938;
#10 a =  4918011965676848001; b =  120488314719630683;
#10 a =  1120294157861489324; b = 5060897469820099834;
#10 a =  8110439193414855071; b =-4655919131134664771;
#10 a =  8158285613393827678; b =-3687499074227118815;
#10 a =  6701463999690318216; b =-2294444897194838689;
#10 a = -8184103843055078809; b =-7165381760252201630;
#10 a =  2014246473658302738; b =-3265716075998056767;
#10 a =  1565875081886578375; b = 2636999868483870953;
#10 a =  6303084787722334955; b = 2679782582529838956;
#10 a =  4556867486542470328; b =-4191124804736556104;
#10 a = -2515157993052333826; b = 7600263886192521676;
#10 a = -3108185468858852085; b = -942424495955610927;
#10 a = -8444393114086798582; b =-5976001838609574441;
#10 a = -8621173582794329215; b =-1718867069814322387;
#10 a =  3180886746062941582; b = 8942354955642713003;
#10 a =  2656307835042104263; b =-5950138324654037501;
#10 a = -7589950408558283838; b =-1642620010659854690;
#10 a = -4513167479626853784; b =-3921971047044787856;
#10 a =  -386264364176222637; b =-1990181519598550773;
#10 a =  4291366351626937070; b =-3099598573668567592;
#10 a =   682399635241269364; b = 2568457296439209466;
#10 a =  3291060271500914736; b =-6484894630511520505;
#10 a = -6218459058794809565; b = 3479470317867366428;
#10 a = -3825962005157280510; b = 7629870895681513356;
#10 a = -3073211819853624231; b = 6297516913852021514;
#10 a =  5406055594701758704; b = 7821451525476900962;
#10 a = -4957614630230187624; b = 8414280879110316540;
#10 a =  7384005035857207052; b =-6004558698365535946;
#10 a =   527598053698037637; b =  560750913630098620;
#10 a =  6934318676579836766; b = -770061046890700591;
#10 a =  8580368801265712150; b =-9154034617326881528;
#10 a =   971414515890299702; b = 3352071459610398210;
#10 a = -2397235868451033504; b =-5838930401611698661;
#10 a =  8733633513794131580; b = 2554780245811100651;
#10 a =  6506951156481937658; b =-5383520875704775974;
#10 a =  -833785339318089305; b =  482375421299610335;
#10 a =  -183276798598995893; b = 6092421285561864235;
#10 a =  5161312971014538908; b =-6756358562559160162;
#10 a =  4143612660497002893; b = 7564334839649471936;
#10 a =  6596549711727760113; b = 3699740822200471067;
#10 a = -7051191807706927123; b =-4191967670633012903;
#10 a =  6094947670178393887; b = 6387802350436752544;
#10 a =  7751058617616963833; b = 5303179114334949532;
#10 a =  9090748793357552486; b =-5591623913352080834;
#10 a =  2955632353434963356; b =-2026947908454003688;
#10 a =  5629927236064746771; b = 3702262460670809808;
#10 a =  8623802675681212330; b = -282854805882528555;
#10 a = -1594012350379521551; b =-8419349307524302221;
#10 a =  4155476075126083224; b =    -942407927874672;
#10 a = -4543419734089236105; b =-7777487071696429114;
#10 a =  8226238535159384540; b =-6697530553640899272;
#10 a = -2923507054760850821; b =-6935874503927689569;
#10 a = -6145717199590563563; b =-7578473078368512650;
#10 a =   718768753143208802; b =-4500722301916392010;
#10 a =   846683107914071167; b =-6305569028175192672;
#10 a = -1874177196043699649; b = 1134744780511356027;
#10 a = -4049740224756722271; b =-4591521175281033345;
#10 a = -9029651167928076594; b =  582462757004215468;
#10 a =  1836743945635871432; b =-6686966105349797094;
#10 a =  3245822879395729737; b =-8055879583975649886;
#10 a = -3817025793818948329; b = 6838456462037737742;
#10 a = -2157121273210247998; b = 8296304405450498645;
#10 a =  1748351954115989507; b = 3304520235116299551;
#10 a =  1161418096130235348; b =-7639482687311991267;
#10 a = -8300891963943693873; b = 7276377954074410654;
#10 a = -8123127662983794232; b =-1322163830127478741;
#10 a = -3478747526507149405; b =-3746897906977754157;
#10 a = -2786679225027643097; b = 7299399861943235082;
#10 a = -7020892249211892690; b =-1212358974979562680;
#10 a =  6100865385405252760; b = 2357047284314947701;
#10 a =  6415998306911286279; b = 2135944322685001663;
#10 a = -2216274628564604961; b =-9039361460003374353;
#10 a =  -195349636612454756; b =-3637088304930198336;
#10 a = -4756070186003321140; b =-1827200295004299727;
#10 a = -5747916621303821512; b = 5399585148706552361;
#10 a =  9138876630020774175; b = 2753449432911047231;
#10 a = -6892161087236908712; b =-7852587821577525704;
#10 a =  1058241618622364700; b = 2134190020689704805;
#10 a =  4834388363920321264; b =-5926451455245703953;
#10 a =  8180895290912051654; b = 1899236512230367930;
#10 a =  9068000165000658357; b =-7702280721760453352;
#10 a = -9162377954293884907; b = 3758199262060734881;
#10 a =  8060059121089389200; b =-6700437061532781062;
#10 a =  6288055369790895076; b = 3330202104324036763;
#10 a = -8547031645487667581; b = 2205498302596829989;
#10 a = -6797707748271016561; b =  997914445667412329;
#10 a =   345031313453332860; b =-3025487350629888352;
#10 a =  3085834908709476451; b = 3347744403309851134;
#10 a =  4810780591521797761; b = 8739201063002623457;
#10 a = -7016380277995124030; b = 5406008028094106637;
#10 a = -2408621924097442865; b = 8349805584016050624;
#10 a = -2483275278490753485; b =-6465057510677709845;
#10 a = -2234845793178346454; b =-1006655144786504966;
#10 a =  2406623827391892756; b =-5050718725059955111;
#10 a = -2098787104809737235; b =-5718877871009420214;
#10 a = -3651848232179750720; b =-8147220605306452285;
#10 a = -2718904862854239299; b = 6498906896546012967;
#10 a =  4700250122219166165; b =-7002231586945497677;
#10 a =   224892719039855821; b =-3248926629264998204;
#10 a = -2472848956102345619; b = 1162445213492607362;
#10 a =  8615091973926745876; b =-5346425258890423556;
#10 a =  3971429073107417323; b = 3119359367511848317;
#10 a = -2635903582352074395; b =-4197739605299044885;
#10 a =   968284810550068923; b =-6970344106666976468;
#10 a =  -397566280808067617; b =  320276304813504544;
#10 a =  6222719457731924551; b =-5443987992787818916;
#10 a =  8996959303770154717; b = 2202535790669742925;
#10 a = -4518538434628558179; b = -753560290115523302;
#10 a = -8981316720151875756; b = 7559516540920142727;
#10 a =  1950674812389868725; b = 8361307801367762848;
#10 a = -1721129064253531821; b =-6369777938184512596;
#10 a = -3625804098905544618; b =-5382983470987149636;
#10 a =  -352937870078893318; b =-8044750659073249471;
#10 a =  6657146787069892874; b =-3770371931435036964;
#10 a = -5117958209645314063; b = 5638565338712617920;
#10 a =  1790946478327042575; b = 4009815765265815049;
#10 a =  2623573435589592786; b =-4063699893818428895;
#10 a =  -288826198686315955; b =-8677249084948046424;
#10 a =   533441427572698758; b =-1050035161663563188;
#10 a =  3159959540599839619; b = 2934952626961057547;
#10 a =   209342588066663696; b = -153604255994961906;
#10 a = -4985554425961020117; b =-4947495010428652066;
#10 a = -4193825429736500083; b =-7926391111558027904;
#10 a = -2323533652716274433; b = 2147598975285705066;
#10 a =   838336616582308408; b =-1760092173766093520;
#10 a =  5273390322895214352; b = 7640210390228003506;
#10 a = -4867643730547242520; b =  415489069122833708;
#10 a = -7720133523843638244; b = 4374239306039125422;
#10 a = -5679095241553023363; b =-8938596440424676585;
#10 a = -3473114208430107074; b =-6554614594105717699;
#10 a = -5433842713593765975; b =-6268582633124258021;
#10 a = -4749827866264157402; b =-5776102415207365630;
#10 a = -2542425478463113766; b = 5509718735691311360;
#10 a =   825643211454431643; b = 7261187850683763122;
#10 a = -1468302767427008423; b = 2877185596176811191;
#10 a =    77466458426838980; b = 7427355452998418433;
#10 a =  7214761631518855020; b = -628908717930043094;
#10 a =  2752119080380880475; b = 5202604719044285369;
#10 a =  5104946191974655643; b =-9056993161546358110;
#10 a =  3398800424525249950; b =-7742521090186675228;
#10 a = -8280768920628764053; b =  782003863996966897;
#10 a = -5757579735000637424; b =-1440444511496051253;
#10 a =  6426851156231796164; b =  555497632592760824;
#10 a =  5356389496433435212; b = 2890910525545030119;
#10 a = -3302397601812713624; b =-5595709790624287679;
#10 a =  2541020333984711106; b = -535734596169881641;
#10 a = -3249142192631932594; b =  743105152333787146;
#10 a =  5132845077250273080; b = 2412510629830672400;
#10 a = -1831784481228827932; b =  292083905101754646;
#10 a =  1247175032471374610; b = 1029983393733845446;
#10 a = -3172189026456945980; b =-7894725379614942912;
#10 a = -8842218448166830244; b = 2864420748528931891;
#10 a =  2288796751368976070; b =-8820374852839363021;
#10 a = -3672552864630790522; b =  638608567159839148;
#10 a =  -546217660709293299; b = 4526218524018067036;
#10 a = -8275410623837294051; b = -314548362085814730;
#10 a = -1053894234665425991; b =-2943098146257508702;
#10 a = -1105083006195194326; b =-5869033999338160357;
#10 a =   -51027553302922749; b = 1202676778649047354;
#10 a = -7312996581380996580; b =-4104925026809896879;
#10 a =   191759815886965563; b =-3406404885814441062;
#10 a = -1414404065311771089; b =-3702248355880983400;
#10 a =  5361951801364729294; b = 7875281243780215014;
#10 a =  7806330156367925995; b =-3136973419043273952;
#10 a = -6095241028324783344; b = 2822027887131234536;
#10 a = -9095017386696782986; b =-1901526427668505526;
#10 a =  8499984743854123202; b =-8692925436407202838;
#10 a = -8246406936366384025; b = 3742541699607072518;
#10 a = -1592644300972322132; b = 8509703077882304616;
#10 a = -7549799940764559970; b = 5417241296288074450;
#10 a =  -830478998237650662; b =-8396017176295884352;
#10 a =  7001211035816942544; b =-8069229967036268050;
#10 a =  8518361870394936115; b = 2962566627123505654;
#10 a = -7912250258896069098; b =-1510760526515615807;
#10 a = -3291118028819853866; b =-5146698104848338939;
#10 a = -5907441254228039330; b =-4691048015157553652;
#10 a =  4017776083546782734; b = 5874138931657612609;
#10 a = -5744076439777312233; b =-3511428239926675115;
#10 a =  8278028390967112152; b = 1690138884875289213;
#10 a =  4241894684584771576; b =-2031555304916776015;
#10 a = -9083158856592762000; b = -994807160166208114;
#10 a = -4299150514137826495; b = 1561756023000781128;
#10 a =  1605153659843328896; b = 8923089418506877685;
#10 a =  5965442865129959054; b =-3745637708034786926;
#10 a = -2481132127946914846; b =-6186459711811479188;
#10 a = -3987388073737486180; b =  -47310517763024454;
#10 a =  2055868983811428878; b =-5437129661355210925;
#10 a =  2270948256434230714; b =  883367512064541310;
#10 a =  6120346650046881371; b =-3908713823064450994;
#10 a = -7541759355763014811; b = 5451859364589988636;
#10 a =   412613155686850161; b =-2663173500824280339;
#10 a =  8982393460914858480; b =-5038207242260564535;
#10 a = -8539381275129743847; b =-3802868961891575893;
#10 a =  7227433061762348724; b = 8960840469624020549;
#10 a = -5905871429810052858; b = 5572255361320382875;
#10 a =  7298000439015835361; b =-1263930950442027698;
#10 a = -4958088341069893208; b = 8217015917502916771;
#10 a =  3469671571612101218; b =-2007004514823644990;
#10 a = -1873091349842506594; b = -258143845702580886;
#10 a = -8108270119505144984; b =-5914908730017353734;
#10 a =  2736726847130018680; b =-8269661611419680654;
#10 a = -1500039205674644625; b =  114945838158034405;
#10 a =  4493267920649267303; b =-5229614891847129769;
#10 a =  8041617476599933419; b = 5656400338486480848;
#10 a =  5221047907427084731; b =-9132738363045073317;
#10 a =  2950777657168263608; b = 1778875774099078144;
#10 a = -8368765064473157925; b = -182774940122464321;
#10 a =   519666694649558817; b =-1464185483970842651;
#10 a =  3656884975470451302; b =-2310342584465107390;
#10 a = -1672738589278186894; b = 2882286022520441881;
#10 a =  -824337824236144962; b = 2805718508073736361;
#10 a =  7703293863662788158; b = 7755474188606652684;
#10 a = -5074737823601292771; b =-5527250211667960358;
#10 a =  9058625699660518660; b = 6236550270475849814;
#10 a = -1207090886735204950; b = 5914159450298426630;
#10 a =  7942848615349404883; b = 9006709560396330841;
#10 a = -3596309370045599339; b = 2291869529673509023;
#10 a =  9212495820271061131; b = 8746140484609937075;
#10 a = -5648951453671261704; b = 8951562527031038150;
#10 a =   107172631289458091; b = -864920298445086098;
#10 a = -2157989791405626465; b =-8194739096879463357;
#10 a =  2197540833410694993; b =-8713847041047459705;
#10 a =  4228870837754928464; b = 8236013276882214124;
#10 a =  8850292333451204597; b = 1047514307267068499;
#10 a = -6294246393611422797; b =-6089193076354782024;
#10 a =  9100517127911213974; b = 4731740845251332208;
#10 a = -7864014048522408092; b = 7331544679458096710;
#10 a = -4153905693968867391; b = 3804024588021470455;
#10 a =  2239490868357687231; b = 5810275572610698972;
#10 a = -3356271628708481565; b =-4042965131472383108;
#10 a =   194573979460193205; b =-3231521574047068912;
#10 a = -3713738735954801687; b =-4565059332955294026;
#10 a =  -697028727988407010; b =-3745920202650043111;
#10 a = -5192243103131210586; b =-1888514347883462468;
#10 a =  8225657571293247393; b =-2186638032012558685;
#10 a = -7032544113453174530; b =-1527772819691394206;
#10 a = -1203197445546142298; b = 4077850855182513987;
#10 a = -7508857328583095320; b = 7239733236149166446;
#10 a = -8018901189445789987; b = 3631735506077857165;
#10 a =  2334820932150086865; b = 5434447514122297233;
#10 a = -2181394218717855242; b = 2204083037587046228;
#10 a =  8700569627852014120; b =-7281808023964204695;
#10 a =   102982341591132423; b = 7038224449669755112;
#10 a =  6232257259655542959; b = 6516455225215342289;
#10 a =  3448924076159565276; b =-2544300127404711313;
#10 a = -6762172233876023992; b =-8088081832152498050;
#10 a =  4687315919463630667; b =-1653726355665356686;
#10 a = -4658369687294119663; b = 6969440785549791775;
#10 a =  1254967729382927147; b = 8823684041337767958;
#10 a =  4833978140635058902; b = 1121532467048439898;
#10 a = -8352498990667805912; b =-3722845922483686525;
#10 a =  4945567939879286640; b =-6632536584944976787;
#10 a = -4832045074451679301; b = 2088867650733565903;
#10 a =  3077989509400455598; b = 5780075913310678801;
#10 a =  6516003823264174344; b =-1952313157950082940;
#10 a = -2954457048260547301; b = -363705043578510228;
#10 a =  1445578430015965204; b =-1347047075453292105;
#10 a =  2792883522389701046; b =-4423396738254726454;
#10 a = -9126000004598227881; b =  -94297809915884363;
#10 a =  8035554086145678624; b = 4630458042348146717;
#10 a =  -216598498611242959; b =-1731892343270218285;
#10 a = -3076825322432085616; b =-8200077805537157991;
#10 a =  5550046711277185365; b =-1410484636833255511;
#10 a = -7094471058877852545; b = 8050918791320235505;
#10 a =  5318593080033274024; b =-4079760893384353008;
#10 a = -6179518653581464676; b = -921180602515140485;
#10 a = -4226855307189332259; b = 8303285674233396027;
#10 a =  3354594208574198689; b = 4192702460709452362;
#10 a =  5466188160894014601; b =-4419626586448574573;
#10 a = -8794359308036076993; b =-4923578970391083196;
#10 a = -8681033922602764745; b =-7068862352871540809;
#10 a = -3842384811408212277; b =-6719193382685102598;
#10 a =  8839802231967662385; b = 7117867216095395754;
#10 a =  3861343176854313171; b = 6613233033935551898;
#10 a = -2224666440069498143; b = 1812662850069117618;
#10 a = -2135185052497565417; b =-8459470301731368717;
#10 a = -8037019423170012092; b = 2753035525738011601;
#10 a = -8626182822230141056; b =-8099873652704512978;
#10 a =   302347921032344884; b =-4553330996911653250;
#10 a =  2824355679280666944; b = 2987525080934473130;
#10 a =  2681777923586821583; b = 3732186579441772083;
#10 a = -3894694240112822505; b =-4520984092174235105;
#10 a =   -45541682473382579; b = -782854773057417467;
#10 a =  6639795317314200348; b = -755175132354670826;
#10 a =   691982178372021386; b = 7757264616208460770;
#10 a =  7530799522014070601; b =-4578505155661293729;
#10 a = -6454349407119862352; b = 7375941960865836125;
#10 a =  5482929734452080381; b =-6025949984396868311;
#10 a =  5823361321139593712; b =-8205684115910581476;
#10 a =  4280580532489573897; b =-6805474626059790533;
#10 a =  3177404798633713760; b = 4215578348360623685;
#10 a =  -604222494886748550; b =  576251962049616845;
#10 a = -8267440842177560062; b =  424436341075076982;
#10 a =  3175012040579255074; b =-7225758947260999111;
#10 a =  1505557930269282400; b =-2895598026137118899;
#10 a =  -166982770860217083; b = 8676226471406281264;
#10 a = -7378749467300822294; b = 4906161565089020293;
#10 a = -6822600187324566912; b = 7889342371621119421;
#10 a =  4274907136413944981; b = 1507260929661647652;
#10 a = -2214053884897213384; b = 8170583454861276208;
#10 a = -4725796690476559400; b = 2969135611088035399;
#10 a =  8316263860220898791; b =-3014338592136057198;
#10 a =  4284892523382830757; b =-1807459522266868752;
#10 a = -1302782155158788690; b =  192396333992311207;
#10 a = -7022401715979190160; b =-3463658440114852185;
#10 a =  5966295235929978613; b =-1095136573795701540;
#10 a = -5872001234569574657; b = -111604197984482815;
#10 a = -2248755758720050032; b = -171772313856205968;
#10 a = -6882952165513303034; b =  276075036519763285;
#10 a = -3909761893188924766; b = 1011509067942964268;
#10 a = -5928253498183157585; b = 6953445346047119162;
#10 a = -6680677227325449295; b =-7056855291162597129;
#10 a =  -110732497011965580; b = 5535418334793347005;
#10 a =  8030308805865963147; b =  858557863670158344;
#10 a =  4713176582910893621; b = 8054320737387908447;
#10 a = -1972334562561986849; b =-3986771122439886849;
#10 a =  7020741068183946638; b = -909317778415806434;
#10 a = -8680589500505928044; b = 7300759988069400423;
#10 a =  7374905641341726164; b = 6114627122346629528;
#10 a = -8977307467630897928; b = 6742985852642927966;
#10 a =  -458939370153904112; b =-8577068242281396091;
#10 a = -5980749831490983391; b =-7604593242072416693;
#10 a =  1719406375501089926; b = 2068543455421053301;
#10 a =  1193380431599843543; b =-5498680729692198208;
#10 a = -2177932476007049868; b =-6473893140009357617;
#10 a =  6256967896733960467; b =-2695997061811609363;
#10 a =   441134814233328884; b = -915857314378017012;
#10 a = -7388038605612941971; b =  163934316778047718;
#10 a = -7383210644626398980; b =-9087294177089479059;
#10 a = -7459683870880179560; b =-5370011227721056053;
#10 a =  6114236316989688825; b = 2833849715446314758;
#10 a =  6210435214893415236; b = 6828551967493249087;
#10 a = -5072500655193616105; b = -440407376238924695;
#10 a =  4172824153155535976; b = 5225380586295990694;
#10 a =   893147053412715824; b =-1394497817599675986;
#10 a =  2897430389442985133; b =-5844060344028082915;
#10 a =  6246496182906832627; b =-1714752736666615777;
#10 a =   258363907008850362; b =-5343067923881493991;
#10 a = -2755054595179788025; b =  669963914226713103;
#10 a = -3220237911566750251; b = 1530680250441555107;
#10 a =  2618243538736035941; b = 1441111373721703936;
    
#10 $finish;
end

initial begin 
    $display( "a,b,sum,carry");
    $monitor( "%d, %d, %d, %b, %b", a, b, sum, cout, OF );
end

initial begin
    $dumpfile( "ripple_carry_64bit.vcd" );
    $dumpvars( 0, RC0 );
end

endmodule